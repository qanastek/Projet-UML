�� {sr  java.io.NotSerializableException(Vx �5  xr java.io.ObjectStreamExceptiond��k�9��  xr java.io.IOExceptionl�sde%�  xr java.lang.Exception��>;�  xr java.lang.Throwable��5'9w�� L causet Ljava/lang/Throwable;L detailMessaget Ljava/lang/String;[ 
stackTracet [Ljava/lang/StackTraceElement;L suppressedExceptionst Ljava/util/List;xpq ~ 	t /src.fr.univavignon.ceri.application.models.Gameur [Ljava.lang.StackTraceElement;F*<<�"9  xp   >sr java.lang.StackTraceElementa	Ś&6݅ I 
lineNumberL declaringClassq ~ L fileNameq ~ L 
methodNameq ~ xp  �t java.io.ObjectOutputStreamt ObjectOutputStream.javat writeObject0sq ~   \q ~ q ~ t writeObjectsq ~   �q ~ 
t 	Game.javat saveGamesq ~    >t 8src.fr.univavignon.ceri.application.EscapeMenuControllert EscapeMenuController.javat savesq ~ ����t $sun.reflect.NativeMethodAccessorImplt NativeMethodAccessorImpl.javat invoke0sq ~    >q ~ q ~ t invokesq ~    +t (sun.reflect.DelegatingMethodAccessorImplt !DelegatingMethodAccessorImpl.javaq ~  sq ~   �t java.lang.reflect.Methodt Method.javaq ~  sq ~    Gt sun.reflect.misc.Trampolinet MethodUtil.javaq ~  sq ~ ����t $sun.reflect.GeneratedMethodAccessor1pq ~  sq ~    +q ~ "q ~ #q ~  sq ~   �q ~ %q ~ &q ~  sq ~   t sun.reflect.misc.MethodUtilq ~ )q ~  sq ~   �t $javafx.fxml.FXMLLoader$MethodHandlert FXMLLoader.javaq ~  sq ~   yt 3javafx.fxml.FXMLLoader$ControllerMethodEventHandlerq ~ 2t handlesq ~    Vt *com.sun.javafx.event.CompositeEventHandlert CompositeEventHandler.javat dispatchBubblingEventsq ~    �t (com.sun.javafx.event.EventHandlerManagert EventHandlerManager.javaq ~ 9sq ~    �q ~ ;q ~ <q ~ 9sq ~    ;t -com.sun.javafx.event.CompositeEventDispatchert CompositeEventDispatcher.javaq ~ 9sq ~    :t )com.sun.javafx.event.BasicEventDispatchert BasicEventDispatcher.javat dispatchEventsq ~    rt +com.sun.javafx.event.EventDispatchChainImplt EventDispatchChainImpl.javaq ~ Dsq ~    8q ~ Bq ~ Cq ~ Dsq ~    rq ~ Fq ~ Gq ~ Dsq ~    8q ~ Bq ~ Cq ~ Dsq ~    rq ~ Fq ~ Gq ~ Dsq ~    Jt com.sun.javafx.event.EventUtilt EventUtil.javat fireEventImplsq ~    1q ~ Mq ~ Nt 	fireEventsq ~    �t javafx.event.Eventt 
Event.javaq ~ Qsq ~    �t javafx.scene.Nodet 	Node.javaq ~ Qsq ~    �t javafx.scene.control.Buttont Button.javat firesq ~    �t 4com.sun.javafx.scene.control.behavior.ButtonBehaviort ButtonBehavior.javat mouseReleasedsq ~    `t 4com.sun.javafx.scene.control.skin.BehaviorSkinBase$1t BehaviorSkinBase.javaq ~ 5sq ~    Yq ~ aq ~ bq ~ 5sq ~    �t Ccom.sun.javafx.event.CompositeEventHandler$NormalEventHandlerRecordq ~ 8t handleBubblingEventsq ~    Pq ~ 7q ~ 8q ~ 9sq ~    �q ~ ;q ~ <q ~ 9sq ~    �q ~ ;q ~ <q ~ 9sq ~    ;q ~ ?q ~ @q ~ 9sq ~    :q ~ Bq ~ Cq ~ Dsq ~    rq ~ Fq ~ Gq ~ Dsq ~    8q ~ Bq ~ Cq ~ Dsq ~    rq ~ Fq ~ Gq ~ Dsq ~    8q ~ Bq ~ Cq ~ Dsq ~    rq ~ Fq ~ Gq ~ Dsq ~    Jq ~ Mq ~ Nq ~ Osq ~    6q ~ Mq ~ Nq ~ Qsq ~    �q ~ Sq ~ Tq ~ Qsq ~   �t javafx.scene.Scene$MouseHandlert 
Scene.javat processsq ~   �q ~ uq ~ vt access$1500sq ~   �t javafx.scene.Sceneq ~ vt impl_processMouseEventsq ~   	�t $javafx.scene.Scene$ScenePeerListenerq ~ vt 
mouseEventsq ~   }t Fcom.sun.javafx.tk.quantum.GlassViewEventHandler$MouseEventNotificationt GlassViewEventHandler.javat runsq ~   'q ~ �q ~ �q ~ �sq ~ ����t java.security.AccessControllert AccessController.javat doPrivilegedsq ~   �t /com.sun.javafx.tk.quantum.GlassViewEventHandlerq ~ �t lambda$handleMouseEvent$354sq ~   �t (com.sun.javafx.tk.quantum.QuantumToolkitt QuantumToolkit.javat runWithoutRenderLocksq ~   �q ~ �q ~ �t handleMouseEventsq ~   +t com.sun.glass.ui.Viewt 	View.javaq ~ �sq ~   �q ~ �q ~ �t notifyMousesq ~ ����t #com.sun.glass.ui.win.WinApplicationt WinApplication.javat _runLoopsq ~    �q ~ �q ~ �t lambda$null$148sq ~   �t java.lang.Threadt Thread.javaq ~ �sr &java.util.Collections$UnmodifiableList�%1�� L listq ~ xr ,java.util.Collections$UnmodifiableCollectionB ��^� L ct Ljava/util/Collection;xpsr java.util.ArrayListx����a� I sizexp    w    xq ~ �x